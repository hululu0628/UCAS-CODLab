`timescale 10ns / 1ns

module custom_cpu(
	input         clk,
	input         rst,

	//Instruction request channel
	output [31:0] PC,
	output        Inst_Req_Valid,
	input         Inst_Req_Ready,

	//Instruction response channel
	input  [31:0] Instruction,
	input         Inst_Valid,
	output        Inst_Ready,

	//Memory request channel
	output [31:0] Address,
	output        MemWrite,
	output [31:0] Write_data,
	output [ 3:0] Write_strb,
	output        MemRead,
	input         Mem_Req_Ready,

	//Memory data response channel
	input  [31:0] Read_data,
	input         Read_data_Valid,
	output        Read_data_Ready,

	input         intr,

	output [31:0] cpu_perf_cnt_0,
	output [31:0] cpu_perf_cnt_1,
	output [31:0] cpu_perf_cnt_2,
	output [31:0] cpu_perf_cnt_3,
	output [31:0] cpu_perf_cnt_4,
	output [31:0] cpu_perf_cnt_5,
	output [31:0] cpu_perf_cnt_6,
	output [31:0] cpu_perf_cnt_7,
	output [31:0] cpu_perf_cnt_8,
	output [31:0] cpu_perf_cnt_9,
	output [31:0] cpu_perf_cnt_10,
	output [31:0] cpu_perf_cnt_11,
	output [31:0] cpu_perf_cnt_12,
	output [31:0] cpu_perf_cnt_13,
	output [31:0] cpu_perf_cnt_14,
	output [31:0] cpu_perf_cnt_15,

	output [69:0] inst_retire
);



/* The following signal is leveraged for behavioral simulation, 
* which is delivered to testbench.
*
* STUDENTS MUST CONTROL LOGICAL BEHAVIORS of THIS SIGNAL.
*
* inst_retired (70-bit): detailed information of the retired instruction,
* mainly including (in order) 
* { 
*   reg_file write-back enable  (69:69,  1-bit),
*   reg_file write-back address (68:64,  5-bit), 
*   reg_file write-back data    (63:32, 32-bit),  
*   retired PC                  (31: 0, 32-bit)
* }
*
*/

	assign inst_retire = {RF_wen,RF_waddr,RF_wdata,PC};//???

  	//wire [69:0] inst_retire;

// TODO: Please add your custom CPU code here
	wire			RF_wen;
	wire [4:0]		RF_waddr;
	wire [31:0]		RF_wdata;

	//divide the instruction into some parts, imm will be generated by instr in Extend
        wire [6:0]opcode;
        wire [4:0]rd,rs1,rs2,shamt;
        wire [2:0]funct3;
        wire [6:0]funct7;
        wire [31:0]inst;
	//determine the type of the instruction
	wire isRtype,isItype_C,isItype_J,isItype_L,isUtype,isJtype,isBtype,isStype;
        wire isShift;
	//change the PC register
	wire PCchange;
	//change the PC register conditionally
	wire PCchangeCond;
	//CU signal
	//without MemWrite and MemRead
	wire RegWrite,MemtoReg,IRWrite,PCWrite,PCWriteCond,ALUsrcA,IorD,PCsrc,Shiftsrc;
	wire [2:0]ALUop,Extype;
	wire [1:0]ALUsrcB;
	
	//some detailed instruction
	wire isbge,isbgeu,isbltu,isblt,isbeq,isbne;
	wire isjalr;
	wire isjal;
	wire islui;
        wire isaulipc;
	//wires using for load instruction
	wire [31:0]W_LoadData,m_MemData;
        wire [31:0]unaligned_Address;
        wire [1:0]offset;
	//wire of register file
	wire [31:0]rdata1,rdata2;
	wire [4:0]raddr1,raddr2;
	//judge if rdata2 = 0
	//should be modified in pipeline
	wire rd1_eq_Zero,rd2_eq_Zero;
	//write_data are selected from these three
	wire [31:0]exwrite,memdatawrite,pcwrite;
	//pc relevant
	wire [31:0]addedpc,nextpc;
	wire PCselect;
        wire [31:0]regPC;

	//store the data fetched from register
	wire [31:0]E_regA,E_regB;

	//the result comes from PC or register file
	wire [31:0]A,B;
	//input of ALU
	//ALU input and output
	wire [2:0]ALUopcode;
	wire [31:0]aluResult;
	wire Overflow,CarryOut,Zero;

	wire [31:0]MW_ExcutionResult,e_ExcutionResult;
	wire W_regZero;

	//decide which op shoule the shifter do
	wire [1:0]Shiftop;
	//shifter input and output
	wire [31:0]shifterA;
	wire [4:0]shifterB;
	wire [31:0]shiftResult;
	//extend output
	wire [31:0]immediate32;

////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


	///*PC Fetch*///
	/*PC register*/
	assign PCchange = PCWrite | PCchangeCond;
	assign PCchangeCond = PCWriteCond & PCselect;
	PC pc(clk,rst,PCchange,nextpc,PC);
        RegisterPC regpc(clk,PC,IRWrite,Inst_Req_Valid,regPC);

	///*Decode*///
	/*Instruction Register*/
	InstructionRegister IR(clk,IRWrite,Instruction,opcode,rd,rs1,rs2,shamt,funct3,funct7,inst);


	assign isRtype = opcode[5] & opcode[4] & ~opcode[2];
	assign isItype_C = ~opcode[5] & opcode[4] & ~opcode[2];
        assign isItype_J = opcode[6] & ~opcode[3] & opcode[2];
        assign isItype_L = ~opcode[5] & ~opcode[4];
        assign isUtype = ~opcode[6] & opcode[2];
        assign isJtype = opcode[3];
        assign isBtype = opcode[6] & ~opcode[2];
        assign isStype = ~opcode[6] & opcode[5] & ~opcode[4];

        assign isShift = ~funct3[1] & funct3[0] & (isRtype | isItype_C);
/*	wire isbge,isbgeu,isbltu,isblt,isbeq,isbne;
	wire isjalr;
	wire isjal;
	wire islui;
        wire isaulipc;
*/
	//instruction
	assign isbge = funct3[2] & ~funct3[1] & funct3[0];
        assign isbgeu = funct3[2] & funct3[1] & funct3[0];
        assign isbltu = funct3[2] & funct3[1] & ~funct3[0];
        assign isblt = funct3[2] & ~funct3[1] & ~funct3[0];
        assign isbeq = ~funct3[2] & ~funct3[1] & ~funct3[0];
        assign isbne = ~funct3[2] & ~funct3[1] & funct3[0];
        assign isjal = isJtype;
        assign isjalr = isItype_J;
        assign isaulipc = ~opcode[6] & ~opcode[5] & opcode[2];
        assign islui = ~opcode[6] & opcode[5] & opcode[2];
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////
	/*Control Unit*/
	ControlUnit control(
	        clk,
	        rst,
	        isRtype,
	        isItype_C,
                isItype_J,
                isItype_L,
                isUtype,
	        isJtype,
	        isBtype,
                isStype, 
                funct3,
                funct7,
	        Inst_Req_Ready,
	        Inst_Valid,
	        Mem_Req_Ready,
	        Read_data_Valid,
	        RegWrite,
	        MemRead,
	        MemWrite,
	        MemtoReg,
	        IRWrite,
	        PCWrite,
	        PCWriteCond,
	        IorD,
	        ALUsrcA,
	        ALUsrcB,
	        Shiftsrc,
	        PCsrc,
                ALUop,
                Extype,
		Inst_Req_Valid,
		Inst_Ready,
		Read_data_Ready,
		cpu_perf_cnt_0,
		cpu_perf_cnt_1,
		cpu_perf_cnt_2,
		cpu_perf_cnt_3,
		cpu_perf_cnt_4,
		cpu_perf_cnt_5,
		cpu_perf_cnt_6,
		cpu_perf_cnt_7,
		cpu_perf_cnt_8
	);
//////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	/*Register File*/
	assign raddr1 = rs1;			//in load and store, rs is base 
	assign raddr2 = rs2;
	//WriteBack
	assign RF_waddr = rd;
	assign memdatawrite = W_LoadData & {32{MemtoReg}};
	assign exwrite = MW_ExcutionResult & {32{~MemtoReg}};
	assign RF_wdata = memdatawrite | exwrite;
	assign RF_wen = RegWrite;

	reg_file register(
		.clk(clk),
		.waddr(RF_waddr),
		.raddr1(raddr1),
		.raddr2(raddr2),
		.wen(RF_wen),
		.wdata(RF_wdata),
		.rdata1(rdata1),
		.rdata2(rdata2)
	);
	RegisterA registerA(clk,rdata1,E_regA);
	RegisterB registerB(clk,rdata2,E_regB);

	///*Excution*///
	/*sign extend*/
	Extend extend(inst,Extype,immediate32);
	/*Shifter*/
	assign Shiftop = {funct7[5],funct3[2]};         //00 is sll,01 is srl,11 is sra
	assign shifterA = E_regA;
	assign shifterB = (E_regB[4:0] & {5{~Shiftsrc}}) | (shamt & {5{Shiftsrc}});
	shifter Shifter(.A(shifterA),.B(shifterB),.Shiftop(Shiftop),.Result(shiftResult));
/////////////////////////////////////////////////////

	/*ALU*/
	//the following two parts are completed in Decoder
	assign A = (E_regA & {32{ALUsrcA}}) | (regPC & {32{~ALUsrcA}});		
	assign B = (E_regB & {32{ALUsrcB[1] & ~ALUsrcB[0]}})
		 | (immediate32 & {32{~ALUsrcB[1]}})
		 | (32'b100 & {32{ALUsrcB[0]}});

	//select a proper operation
	
	alu ALU(.A(A),.B(B),.ALUop(ALUop),.CarryOut(CarryOut),.Overflow(Overflow),.Zero(Zero),.Result(aluResult));

	assign e_ExcutionResult = (aluResult & {32{~islui & ~isShift & ~isItype_J & ~isJtype}}) 
		                | (shiftResult & {32{isShift}})
                                | (immediate32 & {32{islui}})
                                | (PC & {32{isItype_J | isJtype}});
	RegisterALUout aluout(clk,e_ExcutionResult,MW_ExcutionResult);

	
	

	///*MEM*///
	assign Address = ({MW_ExcutionResult[31:2],
                          2'b0} & {32{IorD}}) 
                        | (PC & {32{~IorD}});
        assign offset = MW_ExcutionResult[1:0];
	/*Memory Load*/
	loadData load(.offset(offset),.funct3(funct3),.Read_data(Read_data),.Load_data(m_MemData));
	/*Data Save*/
	storeData store(.offset(offset),.funct3(funct3),.rtdata(rdata2),.Write_data(Write_data),.Write_strb(Write_strb));
	/*MemRegister*/
	RegisterMemData MDR(clk,m_MemData,W_LoadData);



	///*PCupdata*///
	assign addedpc = aluResult;
	//PCsrc & PCWriteCond
	assign PCselect = ((isbeq | isbge | isbgeu) & Zero) | ((isbne | isblt | isbltu) & ~Zero);
	assign nextpc = (MW_ExcutionResult & {32{PCsrc}})
		      | (aluResult & {32{~PCsrc}});


	
endmodule

module PC (
	input clk,
	input rst,
	input PCchange,
	input [31:0]newAddr,
	output reg[31:0]pc
);
	always @(posedge clk)
	begin
		if(rst == 1'b1)
		begin
			pc <= 32'b0;
		end
		else if(PCchange == 1'b1)
		begin
			pc <= newAddr;
		end
		else
			pc <= pc;
	end
endmodule

module Extend(
        input [31:0]inst,
        input [2:0]Extype,
        output [31:0]immediate32
);
	wire imm_31,imm_11,imm_0;
	wire [10:0]imm_30_20;
	wire [7:0]imm_19_12;
	wire [5:0]imm_10_5;
	wire [3:0]imm_4_1;
        wire isIimm,isSimm,isBimm,isUimm,isJimm;

	assign isIimm = ~(|Extype);
        assign isSimm = ~Extype[1] & Extype[0];
        assign isBimm = Extype[1] & ~Extype[0];
        assign isUimm = Extype[2] & ~Extype[0];
        assign isJimm = Extype[1] & Extype[0];

        /*
        assign immI = {{21{inst[31]}},inst[30:25],inst[24:21],inst[20]};
        assign immS = {{21{inst[31]}},inst[30:25],inst[11:8],inst[7]};
        assign immB = {{19{inst[31]}},{2{inst[7]}},inst[30:25],inst[11:8],1'b0};
        assign immU = {inst[31],inst[30:20],inst[19:12],12'b0};
        assign immJ = {{12{inst[31]}},inst[19:12],inst[20],inst[30:25],inst[24:21],1'b0};
        
        

        assign immediate32 = (immI & {32{isIimm}})
                           | (immS & {32{isSimm}})
                           | (immB & {32{isBimm}})
                           | (immU & {32{isUimm}})
                           | (immJ & {32{isJimm}});
	*/
	assign imm_31 = inst[31];
	assign imm_30_20 = {11{inst[31] & ~isUimm}} | (inst[30:20] & {11{isUimm}});
	assign imm_19_12 = {8{inst[31] & ~isUimm & ~isJimm}} | (inst[19:12] & {8{isUimm | isJimm}});
	assign imm_11 = (inst[31] & isIimm) | (inst[31] & isSimm) | (inst[7] & isBimm) | (inst[20] & isJimm);
	assign imm_10_5 = (inst[30:25] & {6{~isUimm}});
	assign imm_4_1 = (inst[24:21] & {4{isIimm | isJimm}}) | (inst[11:8] & {4{isSimm | isBimm}});
	assign imm_0 = (inst[20] & isIimm) | (inst[7] & isSimm);
	assign immediate32 = {imm_31,imm_30_20,imm_19_12,imm_11,imm_10_5,imm_4_1,imm_0};
endmodule
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////
module loadData(
        input [1:0]offset,
	input [2:0]funct3,
	input [31:0]Read_data,
	output [31:0]Load_data
);
	wire [31:0]lb,lh,lw,lbu,lhu;

	//set lb,lh,lw...
        assign lb = {{24{(Read_data[7] & ~offset[1] & ~offset[0]) | (Read_data[15] & ~offset[1] & offset[0])
                        |(Read_data[23] & offset[1] & ~offset[0]) | (Read_data[31] & offset[1] & offset[0])}},
                     ((Read_data[7:0] & {8{~offset[1] & ~offset[0]}}) | (Read_data[15:8] & {8{~offset[1] & offset[0]}})
                     |(Read_data[23:16] & {8{offset[1] & ~offset[0]}}) | (Read_data[31:24] & {8{offset[1] & offset[0]}}))};
        assign lbu = {24'b0,
                      ((Read_data[7:0] & {8{~offset[1] & ~offset[0]}}) | (Read_data[15:8] & {8{~offset[1] & offset[0]}})
                     |(Read_data[23:16] & {8{offset[1] & ~offset[0]}}) | (Read_data[31:24] & {8{offset[1] & offset[0]}}))};
        assign lh = {({16{(Read_data[15] & ~offset[1]) | (Read_data[31] & offset[1])}}),
                     ((Read_data[15:0] & {16{~offset[1]}}) | (Read_data[31:16] & {16{offset[1]}}))};
        assign lhu = {16'b0,((Read_data[15:0] & {16{~offset[1]}}) | (Read_data[31:16] & {16{offset[1]}}))};
        assign lw = Read_data;
	//select the result
        assign Load_data = (lb & {32{~funct3[2] & ~funct3[1] & ~funct3[0]}})
                         | (lbu & {32{funct3[2] & ~funct3[0]}})
                         | (lh & {32{~funct3[2] & funct3[0]}})
                         | (lhu & {32{funct3[2] & funct3[0]}})
                         | (lw & {32{funct3[1]}});
endmodule

module storeData (
        input [1:0]offset,
	input [2:0]funct3,
	input [31:0]rtdata,
	output [31:0]Write_data,
	output [3:0]Write_strb
);
	wire sb,sh,sw;
        wire [31:0]sdata;


        assign sb = ~funct3[1] & ~funct3[0];
        assign sh = funct3[0];
        assign sw = funct3[1];

        assign Write_data = {((rtdata[31:24] & {8{sw}}) | (rtdata[15:8] & {8{sh}}) | (rtdata[7:0] & {8{sb}})),
                             ((rtdata[23:16] & {8{sw}}) | (rtdata[7:0] & {8{sb | sh}})),
                             ((rtdata[15:8] & {8{sw | sh}}) | (rtdata[7:0] & {8{sb}})),
                             (rtdata[7:0])};
        assign Write_strb = {(sw | (sh & offset[1]) | (sb & offset[1] & offset[0])),
                             (sw | (sh & offset[1]) | (sb & offset[1] & ~offset[0])),
                             (sw | (sh & ~offset[1]) | (sb & ~offset[1] & offset[0])),
                             (sw | (sh & ~offset[1]) | (sb & ~offset[1] & ~offset[0]))};

endmodule
////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


module ControlUnit (
	input clk,
	input rst,
	input isRtype,
	input isItype_C,
        input isItype_J,
        input isItype_L,
        input isUtype,
	input isJtype,
	input isBtype,
        input isStype, 
        input [2:0]funct3,
        input [6:0]funct7,
	input Inst_Req_Ready,
	input Inst_Valid,
	input Mem_Req_Ready,
	input Read_data_Valid,
	output RegWrite,
	output MemRead,
	output MemWrite,
	output MemtoReg,
	output IRWrite,
	output PCWrite,
	output PCWriteCond,
	output IorD,
	output ALUsrcA,
	output [1:0]ALUsrcB,
	output Shiftsrc,
	output PCsrc,
        output [2:0]ALUop,
        output [2:0]Extype,
	output Inst_Req_Valid,
	output Inst_Ready,
	output Read_data_Ready,
	output [31:0]cpu_perf_cnt_0,
	output [31:0]cpu_perf_cnt_1,
	output [31:0]cpu_perf_cnt_2,
	output [31:0]cpu_perf_cnt_3,
	output [31:0]cpu_perf_cnt_4,
	output [31:0]cpu_perf_cnt_5,
	output [31:0]cpu_perf_cnt_6,
	output [31:0]cpu_perf_cnt_7,
	output [31:0]cpu_perf_cnt_8
);
	localparam INIT 		= 9'b000000001,	//0
		   IF	 		= 9'b000000010,	//1
		   IW 			= 9'b000000100,	//2
		   ID		 	= 9'b000001000,	//3
		   EX 			= 9'b000010000,	//4
		   ST			= 9'b000100000,	//5
		   LD			= 9'b001000000,	//6
		   RDW			= 9'b010000000,	//7
		   WB			= 9'b100000000;	//8
	
	reg [8:0]current_state,next_state;

	always @(posedge clk)
	begin
		if(rst)
		begin
			current_state <= INIT;
		end
		else
		begin
			current_state <= next_state;
		end
	end

	always @(*)
	begin
		case (current_state)
			INIT:
			begin
				next_state = IF;
			end
			IF:
			begin
				if(Inst_Req_Ready)
					next_state = IW;
				else
					next_state = IF;
				
			end
			IW:
			begin
				if(Inst_Valid)
					next_state = ID;
				else
					next_state = IW;
			end
			ID:
			begin
				next_state = EX;
			end
			EX:
			begin
				if(isRtype | isItype_C | isItype_J | isUtype | isJtype)
					next_state = WB;
				else if(isBtype)
					next_state = IF;
				else if(isStype)
					next_state = ST;
				else if(isItype_L)
					next_state = LD;
				else
					next_state = IF;
			end
			ST:
			begin
				if(Mem_Req_Ready)
					next_state = IF;
				else
					next_state = ST;
			end
			LD:
			begin
				if(Mem_Req_Ready)
					next_state = RDW;
				else
					next_state = LD;
			end
			RDW:
			begin
				if(Read_data_Valid)
					next_state = WB;
				else
					next_state = RDW;
			end
			WB:
			begin
				next_state = IF;
			end
			default: 
				next_state = IF;
		endcase
	end
	/*
	localparam INIT 		= 9'b000000001,	//0
		   IF	 		= 9'b000000010,	//1
		   IW 			= 9'b000000100,	//2
		   ID		 	= 9'b000001000,	//3
		   EX 			= 9'b000010000,	//4
		   ST			= 9'b000100000,	//5
		   LD			= 9'b001000000,	//6
		   RDW			= 9'b010000000,	//7
		   WB			= 9'b100000000;	//8
	*/
	assign IorD 		= current_state[5] | current_state[6];
	assign RegWrite 	= current_state[8] & (isRtype | isUtype | isItype_C | isItype_J | isItype_L | isJtype);
	assign MemRead 		= current_state[6];
	assign MemWrite 	= current_state[5];
	assign MemtoReg 	= current_state[8] & isItype_L;
	assign IRWrite 		= current_state[2] & Inst_Valid;
	assign PCWrite 		= (current_state[4] & (isJtype | isItype_J)) | (current_state[2] & Inst_Valid);
	assign PCWriteCond 	= current_state[4] & (isBtype);
	assign ALUsrcA 		= (|current_state[7:4]) & ~isJtype & ~isUtype;
	assign ALUsrcB 		= (2'b11 & {2{current_state[2]}})
                                | (2'b10 & {2{|current_state[7:4] & (isRtype | isBtype)}});
	assign Shiftsrc 	= isItype_C;
	assign PCsrc 		= current_state[4] & isBtype;
        assign ALUop = (funct3 & {3{(isRtype | isItype_C) & current_state[4]}}) | {2'b0,(isRtype & funct7[5] & current_state[4])}
                     | ({~funct3[2],funct3[2],funct3[1]} & {3{isBtype & current_state[4]}});
        assign Extype           = {isUtype,isBtype,isStype} | {3{isJtype}};
	assign Inst_Req_Valid 	= current_state[1];
	assign Inst_Ready 	= current_state[2] | current_state[0];
	assign Read_data_Ready  = current_state[7] | current_state[0];


	///*Performance Counter*///
	//Runtime cycle count
	reg [31:0] cycle_cnt;
        always @(posedge clk)
        begin
                if(rst)
                        cycle_cnt <= 32'b0;
                else
                        cycle_cnt <= cycle_cnt + 32'b1;
        end
        assign cpu_perf_cnt_0 = cycle_cnt;
	//Instruction count
	reg [31:0] instr_cnt;
	always @(posedge clk)
	begin
		if(rst)
			instr_cnt <= 32'b0;
		else if(current_state[3])
			instr_cnt <= instr_cnt + 32'b1;
		else
			instr_cnt <= instr_cnt;
	end
	assign cpu_perf_cnt_1 = instr_cnt;
	//Instruction request cycle count
	reg [31:0] instr_req_cnt;
	always @(posedge clk)
	begin
		if(rst)
			instr_req_cnt <= 32'b0;
		else if(current_state[1])
			instr_req_cnt <= instr_req_cnt + 32'b1;
		else
			instr_req_cnt <= instr_req_cnt;
	end
	assign cpu_perf_cnt_2 = instr_req_cnt;
	//Instruction valid cycle count
	reg [31:0] instr_valid_cnt;
	always @(posedge clk)
	begin
		if(rst)
			instr_valid_cnt <= 32'b0;
		else if(current_state[2])
			instr_valid_cnt <= instr_valid_cnt + 32'b1;
		else
			instr_valid_cnt <= instr_valid_cnt;
	end
	assign cpu_perf_cnt_3 = instr_valid_cnt;
	//Memory request cycle count(store)
	reg [31:0] mems_req_cnt;
	always @(posedge clk)
	begin
		if(rst)
			mems_req_cnt <= 32'b0;
		else if(current_state[5])
			mems_req_cnt <= mems_req_cnt + 32'b1;
		else
			mems_req_cnt <= mems_req_cnt;
	end
	assign cpu_perf_cnt_4 = mems_req_cnt;
	//Memory request cycle count(load)
	reg [31:0] meml_req_cnt;
	always @(posedge clk)
	begin
		if(rst)
			meml_req_cnt <= 32'b0;
		else if(current_state[6])
			meml_req_cnt <= meml_req_cnt + 32'b1;
		else
			meml_req_cnt <= meml_req_cnt;
	end
	assign cpu_perf_cnt_5 = meml_req_cnt;
	//Memory valid cycle count
	reg [31:0] mem_valid_cnt;
	always @(posedge clk)
	begin
		if(rst)
			mem_valid_cnt <= 32'b0;
		else if(current_state[7])
			mem_valid_cnt <= mem_valid_cnt + 32'b1;
		else
			mem_valid_cnt <= mem_valid_cnt;
	end
	assign cpu_perf_cnt_6 = mem_valid_cnt;
	//Jump count(J-type)
	reg [31:0] jump_cnt;
	always @(posedge clk)
	begin
		if(rst)
			jump_cnt <= 32'b0;
		else if(current_state[4] & (isJtype | isItype_J))
			jump_cnt <= jump_cnt + 32'b1;
		else
			jump_cnt <= jump_cnt;
	end
	assign cpu_perf_cnt_7 = jump_cnt;
	//Branch count(successfully)
	reg [31:0] branch_cnt;
	always @(posedge clk)
	begin
		if(rst)
			branch_cnt <= 32'b0;
		else if(current_state[4] & isBtype)
			branch_cnt <= branch_cnt + 32'b1;
		else
			branch_cnt <= branch_cnt;
	end
	assign cpu_perf_cnt_8 = branch_cnt;

endmodule

module InstructionRegister (
	input clk,
	input IRWrite,
	input [31:0]nextInstruction,
	output [6:0]opcode,
	output [4:0]rd,
	output [4:0]rs1,
	output [4:0]rs2,
	output [4:0]shamt,
	output [2:0]funct3,
        output [6:0]funct7,
        output [31:0]inst
);
	reg [31:0]Instruction;
	always @(posedge clk) begin
		if(IRWrite==1'b1)
			Instruction <= nextInstruction;
		else
			Instruction <= Instruction;
	end

        assign opcode = Instruction[6:0];
        assign rd = Instruction[11:7];
        assign rs1 = Instruction[19:15];
        assign rs2 = Instruction[24:20];
        assign shamt = rs2;
        assign funct3 = Instruction[14:12];
        assign funct7 = Instruction[31:25];
        assign inst = Instruction;

endmodule

module RegisterPC (
        input clk,
        input [31:0]PC,
        input IRWrite,
        input Inst_Req_Valid,
        output [31:0]regPC
);
        reg [31:0]registerpc;
        always @(posedge clk)
        begin
                if(IRWrite == 1'b1 | Inst_Req_Valid==1'b1)
                        registerpc <= PC;
                else
                        registerpc <= registerpc;
        end
        assign regPC = registerpc;
endmodule

module RegisterA (
	input clk,
	input [31:0]rdata1,
	output reg [31:0]E_regA
);
	always @(posedge clk)
	begin
		E_regA <= rdata1;	
	end
	
endmodule

module RegisterB (
	input clk,
	input [31:0]rdata2,
	output reg [31:0]E_regB
);
	always @(posedge clk)
	begin
		E_regB <= rdata2;	
	end
	
endmodule

module RegisterALUout (
	input clk,
	input [31:0]e_ExcutionResult,
	output reg [31:0]MW_ExcutionResult
);
	always @(posedge clk)
	begin
		MW_ExcutionResult <= e_ExcutionResult;	
	end
endmodule

module RegisterZero (
	input clk,
	input Zero,
	output reg W_regZero
);
	always @(posedge clk)
	begin
		W_regZero <= Zero;	
	end
endmodule


module RegisterMemData (
	input clk,
	input [31:0]m_MemData,
	output reg [31:0]W_LoadData
);
	always @(posedge clk)
	begin
		W_LoadData <= m_MemData;	
	end
endmodule
